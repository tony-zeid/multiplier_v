library verilog;
use verilog.vl_types.all;
entity multiplier_v_vlg_vec_tst is
end multiplier_v_vlg_vec_tst;
