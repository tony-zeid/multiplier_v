library verilog;
use verilog.vl_types.all;
entity multiplier_v_vlg_check_tst is
    port(
        pin_name9       : in     vl_logic;
        pin_name10      : in     vl_logic;
        pin_name11      : in     vl_logic;
        pin_name12      : in     vl_logic;
        pin_name13      : in     vl_logic;
        pin_name14      : in     vl_logic;
        pin_name15      : in     vl_logic;
        pin_name16      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end multiplier_v_vlg_check_tst;
