library verilog;
use verilog.vl_types.all;
entity multiplier_v is
    port(
        pin_name9       : out    vl_logic;
        pin_name1       : in     vl_logic;
        pin_name2       : in     vl_logic;
        pin_name3       : in     vl_logic;
        pin_name4       : in     vl_logic;
        pin_name5       : in     vl_logic;
        pin_name6       : in     vl_logic;
        pin_name7       : in     vl_logic;
        pin_name8       : in     vl_logic;
        pin_name10      : out    vl_logic;
        pin_name11      : out    vl_logic;
        pin_name12      : out    vl_logic;
        pin_name13      : out    vl_logic;
        pin_name14      : out    vl_logic;
        pin_name15      : out    vl_logic;
        pin_name16      : out    vl_logic
    );
end multiplier_v;
